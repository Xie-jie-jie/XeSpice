Example ʾ����·
Vin 1 0 10
R1 1 2 1k
R2 2 3 10k
R3 1 3 15k
R4 2 4 40k
R5 3 0 50k
Vmeas 4 0 0
F1 0 3 Vmeas 0.5
.OP
.end

